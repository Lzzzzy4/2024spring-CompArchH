
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h49db1250;
    ram_cell[       1] = 32'h0;  // 32'h86a1c1d9;
    ram_cell[       2] = 32'h0;  // 32'h84922e7a;
    ram_cell[       3] = 32'h0;  // 32'h503f8309;
    ram_cell[       4] = 32'h0;  // 32'he555d029;
    ram_cell[       5] = 32'h0;  // 32'hd73a59a1;
    ram_cell[       6] = 32'h0;  // 32'h83910da4;
    ram_cell[       7] = 32'h0;  // 32'h4180a88e;
    ram_cell[       8] = 32'h0;  // 32'h111ae6bc;
    ram_cell[       9] = 32'h0;  // 32'hcbfe62bf;
    ram_cell[      10] = 32'h0;  // 32'h5b63aa95;
    ram_cell[      11] = 32'h0;  // 32'h46dcc9c6;
    ram_cell[      12] = 32'h0;  // 32'h0844def1;
    ram_cell[      13] = 32'h0;  // 32'h7aaf5234;
    ram_cell[      14] = 32'h0;  // 32'h2a76e8c3;
    ram_cell[      15] = 32'h0;  // 32'h28b2ef56;
    ram_cell[      16] = 32'h0;  // 32'h981cf70b;
    ram_cell[      17] = 32'h0;  // 32'he91d7386;
    ram_cell[      18] = 32'h0;  // 32'hea0e0667;
    ram_cell[      19] = 32'h0;  // 32'hd9b9e28a;
    ram_cell[      20] = 32'h0;  // 32'hbfaa2e8f;
    ram_cell[      21] = 32'h0;  // 32'hdcdbf6c0;
    ram_cell[      22] = 32'h0;  // 32'h1e5485d5;
    ram_cell[      23] = 32'h0;  // 32'h5a31d01d;
    ram_cell[      24] = 32'h0;  // 32'h9866e9d4;
    ram_cell[      25] = 32'h0;  // 32'ha90f7308;
    ram_cell[      26] = 32'h0;  // 32'hf1dbe74d;
    ram_cell[      27] = 32'h0;  // 32'ha026d013;
    ram_cell[      28] = 32'h0;  // 32'hc872ccb1;
    ram_cell[      29] = 32'h0;  // 32'hf71fc9c1;
    ram_cell[      30] = 32'h0;  // 32'h58d588b0;
    ram_cell[      31] = 32'h0;  // 32'h53d55af9;
    ram_cell[      32] = 32'h0;  // 32'h9075cf3a;
    ram_cell[      33] = 32'h0;  // 32'hdaa7c0f6;
    ram_cell[      34] = 32'h0;  // 32'h9bd66920;
    ram_cell[      35] = 32'h0;  // 32'h0eb79772;
    ram_cell[      36] = 32'h0;  // 32'h159864e8;
    ram_cell[      37] = 32'h0;  // 32'h33b61c9d;
    ram_cell[      38] = 32'h0;  // 32'h2947ec5b;
    ram_cell[      39] = 32'h0;  // 32'he60a9f85;
    ram_cell[      40] = 32'h0;  // 32'hf23ea3fd;
    ram_cell[      41] = 32'h0;  // 32'h1ccfc45e;
    ram_cell[      42] = 32'h0;  // 32'h2376d277;
    ram_cell[      43] = 32'h0;  // 32'h57dbf941;
    ram_cell[      44] = 32'h0;  // 32'hf662bbdb;
    ram_cell[      45] = 32'h0;  // 32'ha6b5721f;
    ram_cell[      46] = 32'h0;  // 32'h9f8128cc;
    ram_cell[      47] = 32'h0;  // 32'haa802373;
    ram_cell[      48] = 32'h0;  // 32'h0ba8fd30;
    ram_cell[      49] = 32'h0;  // 32'he302b75e;
    ram_cell[      50] = 32'h0;  // 32'hb56c2b9d;
    ram_cell[      51] = 32'h0;  // 32'h7a445781;
    ram_cell[      52] = 32'h0;  // 32'ha262963f;
    ram_cell[      53] = 32'h0;  // 32'h94c5a5a1;
    ram_cell[      54] = 32'h0;  // 32'he54e10c8;
    ram_cell[      55] = 32'h0;  // 32'hd24b3259;
    ram_cell[      56] = 32'h0;  // 32'hf026b7cb;
    ram_cell[      57] = 32'h0;  // 32'h10abf74a;
    ram_cell[      58] = 32'h0;  // 32'ha298dbba;
    ram_cell[      59] = 32'h0;  // 32'h3f7f0453;
    ram_cell[      60] = 32'h0;  // 32'h02605e08;
    ram_cell[      61] = 32'h0;  // 32'h7f27c408;
    ram_cell[      62] = 32'h0;  // 32'h3ab9b2f9;
    ram_cell[      63] = 32'h0;  // 32'hc7b69d94;
    ram_cell[      64] = 32'h0;  // 32'h5ba696c0;
    ram_cell[      65] = 32'h0;  // 32'hf836adfd;
    ram_cell[      66] = 32'h0;  // 32'h81b0fd8d;
    ram_cell[      67] = 32'h0;  // 32'hf840b679;
    ram_cell[      68] = 32'h0;  // 32'h1b3ea553;
    ram_cell[      69] = 32'h0;  // 32'h2440c1f4;
    ram_cell[      70] = 32'h0;  // 32'hf5c74a1c;
    ram_cell[      71] = 32'h0;  // 32'hb4c79701;
    ram_cell[      72] = 32'h0;  // 32'heee6a9ae;
    ram_cell[      73] = 32'h0;  // 32'h42c1b58e;
    ram_cell[      74] = 32'h0;  // 32'h7bf03bc4;
    ram_cell[      75] = 32'h0;  // 32'h4d043fc5;
    ram_cell[      76] = 32'h0;  // 32'h4f7c2ebd;
    ram_cell[      77] = 32'h0;  // 32'h17de9c27;
    ram_cell[      78] = 32'h0;  // 32'hab5fa3f6;
    ram_cell[      79] = 32'h0;  // 32'h0b36f642;
    ram_cell[      80] = 32'h0;  // 32'h871a2f0c;
    ram_cell[      81] = 32'h0;  // 32'h58d5c3c7;
    ram_cell[      82] = 32'h0;  // 32'h360324ea;
    ram_cell[      83] = 32'h0;  // 32'h6bca1e32;
    ram_cell[      84] = 32'h0;  // 32'he1be5f87;
    ram_cell[      85] = 32'h0;  // 32'h52dee242;
    ram_cell[      86] = 32'h0;  // 32'h6c782f06;
    ram_cell[      87] = 32'h0;  // 32'h22ac7639;
    ram_cell[      88] = 32'h0;  // 32'h2e68c30b;
    ram_cell[      89] = 32'h0;  // 32'h7331a285;
    ram_cell[      90] = 32'h0;  // 32'h8d856f88;
    ram_cell[      91] = 32'h0;  // 32'h7577a871;
    ram_cell[      92] = 32'h0;  // 32'hb82c054c;
    ram_cell[      93] = 32'h0;  // 32'h87823f6c;
    ram_cell[      94] = 32'h0;  // 32'hdd46b803;
    ram_cell[      95] = 32'h0;  // 32'h509db258;
    ram_cell[      96] = 32'h0;  // 32'h438ce04d;
    ram_cell[      97] = 32'h0;  // 32'hcbff4319;
    ram_cell[      98] = 32'h0;  // 32'h8ff5e73f;
    ram_cell[      99] = 32'h0;  // 32'hadd18512;
    ram_cell[     100] = 32'h0;  // 32'h61c46224;
    ram_cell[     101] = 32'h0;  // 32'h4658b068;
    ram_cell[     102] = 32'h0;  // 32'h76765f1b;
    ram_cell[     103] = 32'h0;  // 32'h1b52ee9f;
    ram_cell[     104] = 32'h0;  // 32'hd41db521;
    ram_cell[     105] = 32'h0;  // 32'hfe86001d;
    ram_cell[     106] = 32'h0;  // 32'ha7f618d0;
    ram_cell[     107] = 32'h0;  // 32'hdced7259;
    ram_cell[     108] = 32'h0;  // 32'hb334bd9c;
    ram_cell[     109] = 32'h0;  // 32'h736c2350;
    ram_cell[     110] = 32'h0;  // 32'hd8439735;
    ram_cell[     111] = 32'h0;  // 32'hdc2e5d87;
    ram_cell[     112] = 32'h0;  // 32'h927927e6;
    ram_cell[     113] = 32'h0;  // 32'h36d85903;
    ram_cell[     114] = 32'h0;  // 32'ha15aa5b8;
    ram_cell[     115] = 32'h0;  // 32'habd40e1d;
    ram_cell[     116] = 32'h0;  // 32'hb0efc8dd;
    ram_cell[     117] = 32'h0;  // 32'h7a5f7458;
    ram_cell[     118] = 32'h0;  // 32'h6001655c;
    ram_cell[     119] = 32'h0;  // 32'h2a249411;
    ram_cell[     120] = 32'h0;  // 32'h35383bca;
    ram_cell[     121] = 32'h0;  // 32'h5ceba837;
    ram_cell[     122] = 32'h0;  // 32'h6d51b67d;
    ram_cell[     123] = 32'h0;  // 32'h3ec7fd56;
    ram_cell[     124] = 32'h0;  // 32'h42161c59;
    ram_cell[     125] = 32'h0;  // 32'hf635d5ac;
    ram_cell[     126] = 32'h0;  // 32'h0dfaa556;
    ram_cell[     127] = 32'h0;  // 32'hdd98c1b0;
    ram_cell[     128] = 32'h0;  // 32'h4409620d;
    ram_cell[     129] = 32'h0;  // 32'hb3364742;
    ram_cell[     130] = 32'h0;  // 32'h2d80ddaf;
    ram_cell[     131] = 32'h0;  // 32'h6d4dff4a;
    ram_cell[     132] = 32'h0;  // 32'h73c6303d;
    ram_cell[     133] = 32'h0;  // 32'h5ea59c66;
    ram_cell[     134] = 32'h0;  // 32'h4cdecde3;
    ram_cell[     135] = 32'h0;  // 32'haee91bf7;
    ram_cell[     136] = 32'h0;  // 32'h038af822;
    ram_cell[     137] = 32'h0;  // 32'h3d203a0e;
    ram_cell[     138] = 32'h0;  // 32'h0f4b2dc0;
    ram_cell[     139] = 32'h0;  // 32'h14eaa91e;
    ram_cell[     140] = 32'h0;  // 32'h1cf5d1c0;
    ram_cell[     141] = 32'h0;  // 32'h0908f24a;
    ram_cell[     142] = 32'h0;  // 32'h8cf97c73;
    ram_cell[     143] = 32'h0;  // 32'h897cb7d2;
    ram_cell[     144] = 32'h0;  // 32'hf16358a0;
    ram_cell[     145] = 32'h0;  // 32'ha5be22de;
    ram_cell[     146] = 32'h0;  // 32'hfe52e0a1;
    ram_cell[     147] = 32'h0;  // 32'h642d5ec7;
    ram_cell[     148] = 32'h0;  // 32'h56763cac;
    ram_cell[     149] = 32'h0;  // 32'h2b2cade1;
    ram_cell[     150] = 32'h0;  // 32'h93c4e2b0;
    ram_cell[     151] = 32'h0;  // 32'h6281d5d9;
    ram_cell[     152] = 32'h0;  // 32'hb1bb15d3;
    ram_cell[     153] = 32'h0;  // 32'hadcc967d;
    ram_cell[     154] = 32'h0;  // 32'h9ee1651c;
    ram_cell[     155] = 32'h0;  // 32'h9223f741;
    ram_cell[     156] = 32'h0;  // 32'hfd7f4aee;
    ram_cell[     157] = 32'h0;  // 32'h44158503;
    ram_cell[     158] = 32'h0;  // 32'h91be5746;
    ram_cell[     159] = 32'h0;  // 32'hcdf3bdac;
    ram_cell[     160] = 32'h0;  // 32'h96e2c51d;
    ram_cell[     161] = 32'h0;  // 32'h284f03a5;
    ram_cell[     162] = 32'h0;  // 32'h858d9c38;
    ram_cell[     163] = 32'h0;  // 32'hc29523b2;
    ram_cell[     164] = 32'h0;  // 32'ha9cf0503;
    ram_cell[     165] = 32'h0;  // 32'h2999d8da;
    ram_cell[     166] = 32'h0;  // 32'h35ab017e;
    ram_cell[     167] = 32'h0;  // 32'h5a515640;
    ram_cell[     168] = 32'h0;  // 32'he7ff0f52;
    ram_cell[     169] = 32'h0;  // 32'h25b860ae;
    ram_cell[     170] = 32'h0;  // 32'h5733817a;
    ram_cell[     171] = 32'h0;  // 32'haa878649;
    ram_cell[     172] = 32'h0;  // 32'h3f4cbb2d;
    ram_cell[     173] = 32'h0;  // 32'h4381f165;
    ram_cell[     174] = 32'h0;  // 32'hf7148bfc;
    ram_cell[     175] = 32'h0;  // 32'hf0553b08;
    ram_cell[     176] = 32'h0;  // 32'h747257a9;
    ram_cell[     177] = 32'h0;  // 32'hfea9b827;
    ram_cell[     178] = 32'h0;  // 32'h7f2f10ef;
    ram_cell[     179] = 32'h0;  // 32'he0b7ca9b;
    ram_cell[     180] = 32'h0;  // 32'h67ad59df;
    ram_cell[     181] = 32'h0;  // 32'h571e66c4;
    ram_cell[     182] = 32'h0;  // 32'h6027868a;
    ram_cell[     183] = 32'h0;  // 32'h39bc719e;
    ram_cell[     184] = 32'h0;  // 32'h2beaaa60;
    ram_cell[     185] = 32'h0;  // 32'h188616a3;
    ram_cell[     186] = 32'h0;  // 32'h786cf1b4;
    ram_cell[     187] = 32'h0;  // 32'h3cfdc84b;
    ram_cell[     188] = 32'h0;  // 32'heb25a852;
    ram_cell[     189] = 32'h0;  // 32'hb098a860;
    ram_cell[     190] = 32'h0;  // 32'h36364496;
    ram_cell[     191] = 32'h0;  // 32'h13f969fe;
    ram_cell[     192] = 32'h0;  // 32'hd292954b;
    ram_cell[     193] = 32'h0;  // 32'h911518a5;
    ram_cell[     194] = 32'h0;  // 32'he6dfbbf1;
    ram_cell[     195] = 32'h0;  // 32'hb488eb7a;
    ram_cell[     196] = 32'h0;  // 32'ha0342472;
    ram_cell[     197] = 32'h0;  // 32'h57091b61;
    ram_cell[     198] = 32'h0;  // 32'hfc59c707;
    ram_cell[     199] = 32'h0;  // 32'h0a566869;
    ram_cell[     200] = 32'h0;  // 32'ha0e783c7;
    ram_cell[     201] = 32'h0;  // 32'h4620025d;
    ram_cell[     202] = 32'h0;  // 32'hfe01d7df;
    ram_cell[     203] = 32'h0;  // 32'h42d89112;
    ram_cell[     204] = 32'h0;  // 32'h8a23bac0;
    ram_cell[     205] = 32'h0;  // 32'ha69f8786;
    ram_cell[     206] = 32'h0;  // 32'h9b1d6fc2;
    ram_cell[     207] = 32'h0;  // 32'h2ae2b0e5;
    ram_cell[     208] = 32'h0;  // 32'h3df6632a;
    ram_cell[     209] = 32'h0;  // 32'h7683714a;
    ram_cell[     210] = 32'h0;  // 32'h23ea13a1;
    ram_cell[     211] = 32'h0;  // 32'h0aa7c54b;
    ram_cell[     212] = 32'h0;  // 32'h75a0afaa;
    ram_cell[     213] = 32'h0;  // 32'h4fb1745c;
    ram_cell[     214] = 32'h0;  // 32'hecf43aed;
    ram_cell[     215] = 32'h0;  // 32'h4527666d;
    ram_cell[     216] = 32'h0;  // 32'h6c00dc76;
    ram_cell[     217] = 32'h0;  // 32'h519d46db;
    ram_cell[     218] = 32'h0;  // 32'hbe9de764;
    ram_cell[     219] = 32'h0;  // 32'hd0361d96;
    ram_cell[     220] = 32'h0;  // 32'h2a145dea;
    ram_cell[     221] = 32'h0;  // 32'h974385f7;
    ram_cell[     222] = 32'h0;  // 32'h4dcc3a11;
    ram_cell[     223] = 32'h0;  // 32'he65f69fc;
    ram_cell[     224] = 32'h0;  // 32'h7bfdeb49;
    ram_cell[     225] = 32'h0;  // 32'he97fd79f;
    ram_cell[     226] = 32'h0;  // 32'h4a8e13a4;
    ram_cell[     227] = 32'h0;  // 32'h4c0e4878;
    ram_cell[     228] = 32'h0;  // 32'h00f379fa;
    ram_cell[     229] = 32'h0;  // 32'he9191b4a;
    ram_cell[     230] = 32'h0;  // 32'h557f46f1;
    ram_cell[     231] = 32'h0;  // 32'h435e7a77;
    ram_cell[     232] = 32'h0;  // 32'he884bddb;
    ram_cell[     233] = 32'h0;  // 32'hb5784437;
    ram_cell[     234] = 32'h0;  // 32'h748b1df7;
    ram_cell[     235] = 32'h0;  // 32'h8b660bca;
    ram_cell[     236] = 32'h0;  // 32'h31d150d3;
    ram_cell[     237] = 32'h0;  // 32'hcc8466cb;
    ram_cell[     238] = 32'h0;  // 32'hb8da3ac0;
    ram_cell[     239] = 32'h0;  // 32'hddb37098;
    ram_cell[     240] = 32'h0;  // 32'hcd6683c8;
    ram_cell[     241] = 32'h0;  // 32'h3afb00aa;
    ram_cell[     242] = 32'h0;  // 32'hbc8eec39;
    ram_cell[     243] = 32'h0;  // 32'hfca16c2d;
    ram_cell[     244] = 32'h0;  // 32'hf83e744e;
    ram_cell[     245] = 32'h0;  // 32'ha3bc73af;
    ram_cell[     246] = 32'h0;  // 32'hf237e4c6;
    ram_cell[     247] = 32'h0;  // 32'h87387a25;
    ram_cell[     248] = 32'h0;  // 32'h51483163;
    ram_cell[     249] = 32'h0;  // 32'h6aa04e1a;
    ram_cell[     250] = 32'h0;  // 32'h5dd16776;
    ram_cell[     251] = 32'h0;  // 32'h28b352aa;
    ram_cell[     252] = 32'h0;  // 32'h1672f417;
    ram_cell[     253] = 32'h0;  // 32'h82b09cd4;
    ram_cell[     254] = 32'h0;  // 32'hafc279a9;
    ram_cell[     255] = 32'h0;  // 32'hbf47269b;
    // src matrix A
    ram_cell[     256] = 32'h044c0c9a;
    ram_cell[     257] = 32'h38461078;
    ram_cell[     258] = 32'haf38ef4c;
    ram_cell[     259] = 32'h052b614c;
    ram_cell[     260] = 32'h296056f0;
    ram_cell[     261] = 32'h67efbccd;
    ram_cell[     262] = 32'h52e88c5b;
    ram_cell[     263] = 32'h53186079;
    ram_cell[     264] = 32'h7936cacd;
    ram_cell[     265] = 32'h8ff98a8c;
    ram_cell[     266] = 32'hefb53232;
    ram_cell[     267] = 32'hdbad2bf2;
    ram_cell[     268] = 32'h455e4755;
    ram_cell[     269] = 32'ha39a2df3;
    ram_cell[     270] = 32'h2ea67600;
    ram_cell[     271] = 32'h8377f03b;
    ram_cell[     272] = 32'hd9b822de;
    ram_cell[     273] = 32'h3b211484;
    ram_cell[     274] = 32'h9593e80d;
    ram_cell[     275] = 32'h0d56f4c6;
    ram_cell[     276] = 32'h3cbd0ddf;
    ram_cell[     277] = 32'hc54d9fd4;
    ram_cell[     278] = 32'hc58ae42e;
    ram_cell[     279] = 32'h7f6baafd;
    ram_cell[     280] = 32'hf67245f2;
    ram_cell[     281] = 32'h67c935b0;
    ram_cell[     282] = 32'h747e5b64;
    ram_cell[     283] = 32'h27f0349e;
    ram_cell[     284] = 32'h4e21a008;
    ram_cell[     285] = 32'h6c59d95c;
    ram_cell[     286] = 32'h9f9b0130;
    ram_cell[     287] = 32'h9195ac99;
    ram_cell[     288] = 32'hfc36a65a;
    ram_cell[     289] = 32'h97f19c55;
    ram_cell[     290] = 32'h46180c86;
    ram_cell[     291] = 32'h097fe8cd;
    ram_cell[     292] = 32'h70748447;
    ram_cell[     293] = 32'h3304a8dd;
    ram_cell[     294] = 32'h8f8dde1b;
    ram_cell[     295] = 32'h73990b1d;
    ram_cell[     296] = 32'h3f947ddc;
    ram_cell[     297] = 32'h2de7df03;
    ram_cell[     298] = 32'hf2f51140;
    ram_cell[     299] = 32'h5d0d4b3b;
    ram_cell[     300] = 32'h80821349;
    ram_cell[     301] = 32'had798f27;
    ram_cell[     302] = 32'h793e136e;
    ram_cell[     303] = 32'hcb9a7c49;
    ram_cell[     304] = 32'h2c471d5c;
    ram_cell[     305] = 32'hf0d6d60b;
    ram_cell[     306] = 32'hed1dd488;
    ram_cell[     307] = 32'hc29fe40b;
    ram_cell[     308] = 32'h50b2e682;
    ram_cell[     309] = 32'h2bd6b3b5;
    ram_cell[     310] = 32'hff4b2f65;
    ram_cell[     311] = 32'ha0a03663;
    ram_cell[     312] = 32'h8eeb4c6f;
    ram_cell[     313] = 32'h76f6c905;
    ram_cell[     314] = 32'ha38ff9b4;
    ram_cell[     315] = 32'hf0990728;
    ram_cell[     316] = 32'h8a9b206b;
    ram_cell[     317] = 32'hec1f5585;
    ram_cell[     318] = 32'h8126faa6;
    ram_cell[     319] = 32'hfdc91288;
    ram_cell[     320] = 32'he2fb2c06;
    ram_cell[     321] = 32'hb3588504;
    ram_cell[     322] = 32'hf4efba8f;
    ram_cell[     323] = 32'hb6c74e72;
    ram_cell[     324] = 32'h3bab8d72;
    ram_cell[     325] = 32'hbd26427c;
    ram_cell[     326] = 32'ha7f5befc;
    ram_cell[     327] = 32'hd3368eed;
    ram_cell[     328] = 32'h3c5f97e0;
    ram_cell[     329] = 32'h75cc0958;
    ram_cell[     330] = 32'h94ed074b;
    ram_cell[     331] = 32'h1c15fc64;
    ram_cell[     332] = 32'h48f3655d;
    ram_cell[     333] = 32'hea3750ce;
    ram_cell[     334] = 32'h0ac51d8b;
    ram_cell[     335] = 32'hdd6c4bbd;
    ram_cell[     336] = 32'h63ec8b10;
    ram_cell[     337] = 32'hb8d3253b;
    ram_cell[     338] = 32'h0eb715c2;
    ram_cell[     339] = 32'hc1df8241;
    ram_cell[     340] = 32'h30e89718;
    ram_cell[     341] = 32'h1eb6e310;
    ram_cell[     342] = 32'hb3467957;
    ram_cell[     343] = 32'hb185291f;
    ram_cell[     344] = 32'hc3462267;
    ram_cell[     345] = 32'hd72a84e3;
    ram_cell[     346] = 32'h46579197;
    ram_cell[     347] = 32'h0576e9d5;
    ram_cell[     348] = 32'h19c9cf51;
    ram_cell[     349] = 32'h0bc41348;
    ram_cell[     350] = 32'ha8d8b470;
    ram_cell[     351] = 32'h7541db46;
    ram_cell[     352] = 32'h691b2975;
    ram_cell[     353] = 32'h9331d44d;
    ram_cell[     354] = 32'h05d2d1cb;
    ram_cell[     355] = 32'h2f0092aa;
    ram_cell[     356] = 32'h9e207212;
    ram_cell[     357] = 32'hf0499b69;
    ram_cell[     358] = 32'h3c5df60c;
    ram_cell[     359] = 32'h4bdd2cf2;
    ram_cell[     360] = 32'h47be2c1a;
    ram_cell[     361] = 32'hf7fc204f;
    ram_cell[     362] = 32'hccf86a75;
    ram_cell[     363] = 32'hb077c6a7;
    ram_cell[     364] = 32'h224c6713;
    ram_cell[     365] = 32'h161b8c63;
    ram_cell[     366] = 32'h5029364d;
    ram_cell[     367] = 32'ha8c8258d;
    ram_cell[     368] = 32'h5883bff9;
    ram_cell[     369] = 32'h62beeb08;
    ram_cell[     370] = 32'h55e6b683;
    ram_cell[     371] = 32'h9c7266fc;
    ram_cell[     372] = 32'h818d9b87;
    ram_cell[     373] = 32'h703d2401;
    ram_cell[     374] = 32'h1aa8e2c5;
    ram_cell[     375] = 32'h02907008;
    ram_cell[     376] = 32'h87f143fa;
    ram_cell[     377] = 32'hc402407a;
    ram_cell[     378] = 32'h67719050;
    ram_cell[     379] = 32'h8c2b6db1;
    ram_cell[     380] = 32'hf97c4421;
    ram_cell[     381] = 32'hb8f03160;
    ram_cell[     382] = 32'hb3954430;
    ram_cell[     383] = 32'h3dde21ee;
    ram_cell[     384] = 32'h282965f3;
    ram_cell[     385] = 32'heaf96cd5;
    ram_cell[     386] = 32'hf69aa596;
    ram_cell[     387] = 32'hd242428d;
    ram_cell[     388] = 32'h355e2811;
    ram_cell[     389] = 32'h3e2c379b;
    ram_cell[     390] = 32'hf687867d;
    ram_cell[     391] = 32'he67fd641;
    ram_cell[     392] = 32'hf08d989a;
    ram_cell[     393] = 32'he8cae990;
    ram_cell[     394] = 32'h4cf9b431;
    ram_cell[     395] = 32'h0ebeecf4;
    ram_cell[     396] = 32'h53b622f5;
    ram_cell[     397] = 32'h4569249a;
    ram_cell[     398] = 32'h6acb542b;
    ram_cell[     399] = 32'h9e63b3ce;
    ram_cell[     400] = 32'h22f8ecc4;
    ram_cell[     401] = 32'h035481e1;
    ram_cell[     402] = 32'h93d7f0d5;
    ram_cell[     403] = 32'h5983d3e3;
    ram_cell[     404] = 32'hfdad6f98;
    ram_cell[     405] = 32'hc3af396e;
    ram_cell[     406] = 32'hd5aab528;
    ram_cell[     407] = 32'h75363c84;
    ram_cell[     408] = 32'h1fcba071;
    ram_cell[     409] = 32'h315c7033;
    ram_cell[     410] = 32'ha2f0a7c5;
    ram_cell[     411] = 32'hec76a5d5;
    ram_cell[     412] = 32'hc884e738;
    ram_cell[     413] = 32'h977a2d76;
    ram_cell[     414] = 32'h9ce2dc0c;
    ram_cell[     415] = 32'h59fdf08b;
    ram_cell[     416] = 32'h51f9f582;
    ram_cell[     417] = 32'h15f4fa6f;
    ram_cell[     418] = 32'h6a838089;
    ram_cell[     419] = 32'h6a6626be;
    ram_cell[     420] = 32'hfb2aa9c3;
    ram_cell[     421] = 32'hcb38567f;
    ram_cell[     422] = 32'ha245b0d5;
    ram_cell[     423] = 32'h4dcc3d8f;
    ram_cell[     424] = 32'hba57546a;
    ram_cell[     425] = 32'h2a087a5b;
    ram_cell[     426] = 32'h171c53d0;
    ram_cell[     427] = 32'h7a0e58c4;
    ram_cell[     428] = 32'h85381e9e;
    ram_cell[     429] = 32'h16376447;
    ram_cell[     430] = 32'he1afa65d;
    ram_cell[     431] = 32'h888e9082;
    ram_cell[     432] = 32'h386ab53a;
    ram_cell[     433] = 32'h6ccda62d;
    ram_cell[     434] = 32'hdcab0644;
    ram_cell[     435] = 32'h1010473e;
    ram_cell[     436] = 32'h038e0bd3;
    ram_cell[     437] = 32'h50957cff;
    ram_cell[     438] = 32'h577aa071;
    ram_cell[     439] = 32'h81117cd5;
    ram_cell[     440] = 32'ha68b7f49;
    ram_cell[     441] = 32'h7163d63c;
    ram_cell[     442] = 32'h3419d35d;
    ram_cell[     443] = 32'he4bc37c9;
    ram_cell[     444] = 32'h7ff89da0;
    ram_cell[     445] = 32'h1b8c7383;
    ram_cell[     446] = 32'hc488923c;
    ram_cell[     447] = 32'h77170bef;
    ram_cell[     448] = 32'h9f096dc0;
    ram_cell[     449] = 32'h849fb2c8;
    ram_cell[     450] = 32'h24e6e478;
    ram_cell[     451] = 32'hd2925662;
    ram_cell[     452] = 32'hc5e18e5e;
    ram_cell[     453] = 32'h51685457;
    ram_cell[     454] = 32'he0e5161c;
    ram_cell[     455] = 32'ha2121bf7;
    ram_cell[     456] = 32'h672d1867;
    ram_cell[     457] = 32'h89057c5d;
    ram_cell[     458] = 32'hbb6842b8;
    ram_cell[     459] = 32'h9c6f99e3;
    ram_cell[     460] = 32'hcbe0c526;
    ram_cell[     461] = 32'h123d262d;
    ram_cell[     462] = 32'hd7c9f1cf;
    ram_cell[     463] = 32'hf6d4818f;
    ram_cell[     464] = 32'h66c8faef;
    ram_cell[     465] = 32'h0c2a8cfb;
    ram_cell[     466] = 32'hfa7a1a69;
    ram_cell[     467] = 32'hb8e54512;
    ram_cell[     468] = 32'had78702c;
    ram_cell[     469] = 32'h15f6990f;
    ram_cell[     470] = 32'hcfd40a96;
    ram_cell[     471] = 32'h57c01fe4;
    ram_cell[     472] = 32'h99cde6f1;
    ram_cell[     473] = 32'h796e05f1;
    ram_cell[     474] = 32'he4786720;
    ram_cell[     475] = 32'hd059a6b8;
    ram_cell[     476] = 32'hef7cda8a;
    ram_cell[     477] = 32'h5f9328e1;
    ram_cell[     478] = 32'h4e61d6fa;
    ram_cell[     479] = 32'h4bbb4f0d;
    ram_cell[     480] = 32'hd7dab1b3;
    ram_cell[     481] = 32'h60c9535f;
    ram_cell[     482] = 32'hc3d17acd;
    ram_cell[     483] = 32'h9c99e901;
    ram_cell[     484] = 32'h7607f80d;
    ram_cell[     485] = 32'hee90f287;
    ram_cell[     486] = 32'hc19ca4bd;
    ram_cell[     487] = 32'hf02a205b;
    ram_cell[     488] = 32'hf7971261;
    ram_cell[     489] = 32'hb3458d38;
    ram_cell[     490] = 32'h50dee9d2;
    ram_cell[     491] = 32'h037fc92d;
    ram_cell[     492] = 32'h4d363c72;
    ram_cell[     493] = 32'h54d47204;
    ram_cell[     494] = 32'ha5dfc2ec;
    ram_cell[     495] = 32'h4b417906;
    ram_cell[     496] = 32'hc677da0d;
    ram_cell[     497] = 32'h68fb2f84;
    ram_cell[     498] = 32'hb786576c;
    ram_cell[     499] = 32'h81b1134f;
    ram_cell[     500] = 32'h4a470e23;
    ram_cell[     501] = 32'h07c6cb4c;
    ram_cell[     502] = 32'h02670c2e;
    ram_cell[     503] = 32'hb9e5d371;
    ram_cell[     504] = 32'h6a11862c;
    ram_cell[     505] = 32'h877c365e;
    ram_cell[     506] = 32'h076cf4d9;
    ram_cell[     507] = 32'h9b7d3630;
    ram_cell[     508] = 32'h40edbf82;
    ram_cell[     509] = 32'h037a3ae0;
    ram_cell[     510] = 32'hd7273dd2;
    ram_cell[     511] = 32'h8f6f2981;
    // src matrix B
    ram_cell[     512] = 32'h6e2e702f;
    ram_cell[     513] = 32'h2db13936;
    ram_cell[     514] = 32'h3a4b27d8;
    ram_cell[     515] = 32'h5301a610;
    ram_cell[     516] = 32'he6053c29;
    ram_cell[     517] = 32'hed378ea4;
    ram_cell[     518] = 32'h71bb383f;
    ram_cell[     519] = 32'hf27e64a7;
    ram_cell[     520] = 32'h0dba7eb7;
    ram_cell[     521] = 32'hf13b54e3;
    ram_cell[     522] = 32'h28dcb475;
    ram_cell[     523] = 32'ha1724b90;
    ram_cell[     524] = 32'hcbc85ee4;
    ram_cell[     525] = 32'h987e308b;
    ram_cell[     526] = 32'hb8569b79;
    ram_cell[     527] = 32'hbac91eba;
    ram_cell[     528] = 32'h2d26f41e;
    ram_cell[     529] = 32'h0a856a34;
    ram_cell[     530] = 32'h30e93a2b;
    ram_cell[     531] = 32'hb8dbc0c5;
    ram_cell[     532] = 32'hd21c4cca;
    ram_cell[     533] = 32'h3f538aef;
    ram_cell[     534] = 32'h62eb3551;
    ram_cell[     535] = 32'h512dca22;
    ram_cell[     536] = 32'h93fd1d4b;
    ram_cell[     537] = 32'h1c6ed551;
    ram_cell[     538] = 32'h8e29f488;
    ram_cell[     539] = 32'h71bc1d95;
    ram_cell[     540] = 32'ha85550bb;
    ram_cell[     541] = 32'h0b10e1a3;
    ram_cell[     542] = 32'h8787e9d6;
    ram_cell[     543] = 32'hf5bf857b;
    ram_cell[     544] = 32'hcd5ab6c7;
    ram_cell[     545] = 32'h0b1cc32c;
    ram_cell[     546] = 32'hf9fc2409;
    ram_cell[     547] = 32'h86142809;
    ram_cell[     548] = 32'h66c55d37;
    ram_cell[     549] = 32'hef451aae;
    ram_cell[     550] = 32'h2da9e7da;
    ram_cell[     551] = 32'h3448ec94;
    ram_cell[     552] = 32'hed48f51e;
    ram_cell[     553] = 32'hbfab1d07;
    ram_cell[     554] = 32'h58a5775d;
    ram_cell[     555] = 32'hf3b25dc3;
    ram_cell[     556] = 32'hc268e9b3;
    ram_cell[     557] = 32'hb5a028f0;
    ram_cell[     558] = 32'hf5982fed;
    ram_cell[     559] = 32'hf5ffb2b7;
    ram_cell[     560] = 32'heed84517;
    ram_cell[     561] = 32'h1415ba2b;
    ram_cell[     562] = 32'hfe3f7ff3;
    ram_cell[     563] = 32'h6736f435;
    ram_cell[     564] = 32'h4f6540eb;
    ram_cell[     565] = 32'he57944c0;
    ram_cell[     566] = 32'h3c93a810;
    ram_cell[     567] = 32'h90f0e2f9;
    ram_cell[     568] = 32'h7a8ae258;
    ram_cell[     569] = 32'hc6f9c26e;
    ram_cell[     570] = 32'h1cece573;
    ram_cell[     571] = 32'h1cdfcb8d;
    ram_cell[     572] = 32'hbadd7d7c;
    ram_cell[     573] = 32'hd8fb685b;
    ram_cell[     574] = 32'hb501ff14;
    ram_cell[     575] = 32'h018100e2;
    ram_cell[     576] = 32'h5ac91f9b;
    ram_cell[     577] = 32'hd8aaefbe;
    ram_cell[     578] = 32'hd73934bb;
    ram_cell[     579] = 32'h6bd8e38d;
    ram_cell[     580] = 32'h38d89f37;
    ram_cell[     581] = 32'h5d2ddfe6;
    ram_cell[     582] = 32'hf8b0568b;
    ram_cell[     583] = 32'haddcfa12;
    ram_cell[     584] = 32'hebc9afd1;
    ram_cell[     585] = 32'h944e1713;
    ram_cell[     586] = 32'h0ed5fe17;
    ram_cell[     587] = 32'h8c3cf045;
    ram_cell[     588] = 32'h719dbe01;
    ram_cell[     589] = 32'h07dd3a45;
    ram_cell[     590] = 32'ha64a69b2;
    ram_cell[     591] = 32'h6f458be0;
    ram_cell[     592] = 32'h1fad5768;
    ram_cell[     593] = 32'h87cf0620;
    ram_cell[     594] = 32'hfb0dfaf3;
    ram_cell[     595] = 32'hfa30495b;
    ram_cell[     596] = 32'h129606a0;
    ram_cell[     597] = 32'h53f6946f;
    ram_cell[     598] = 32'h5c11068d;
    ram_cell[     599] = 32'h893e3d95;
    ram_cell[     600] = 32'h3acc89de;
    ram_cell[     601] = 32'he1c6deb3;
    ram_cell[     602] = 32'h281b2541;
    ram_cell[     603] = 32'h9c90ea8f;
    ram_cell[     604] = 32'h2d60293b;
    ram_cell[     605] = 32'h6d7d4a12;
    ram_cell[     606] = 32'hfa31ba3a;
    ram_cell[     607] = 32'h76280585;
    ram_cell[     608] = 32'ha14042a5;
    ram_cell[     609] = 32'haaa9881e;
    ram_cell[     610] = 32'he3288568;
    ram_cell[     611] = 32'h28b8251b;
    ram_cell[     612] = 32'hd2cd6591;
    ram_cell[     613] = 32'hb695cc26;
    ram_cell[     614] = 32'hc2236deb;
    ram_cell[     615] = 32'hd3dc5ed7;
    ram_cell[     616] = 32'h57e892ce;
    ram_cell[     617] = 32'h3881a911;
    ram_cell[     618] = 32'hb2363389;
    ram_cell[     619] = 32'hf0feddd9;
    ram_cell[     620] = 32'h7deef036;
    ram_cell[     621] = 32'he2460beb;
    ram_cell[     622] = 32'h1e51b5ec;
    ram_cell[     623] = 32'ha8880268;
    ram_cell[     624] = 32'h56cb44b5;
    ram_cell[     625] = 32'h8cdebc8c;
    ram_cell[     626] = 32'hc07a15ee;
    ram_cell[     627] = 32'h0b0cdad7;
    ram_cell[     628] = 32'hfb2a9a94;
    ram_cell[     629] = 32'h4d9bc270;
    ram_cell[     630] = 32'h099761ac;
    ram_cell[     631] = 32'h526728f1;
    ram_cell[     632] = 32'h9d7a401a;
    ram_cell[     633] = 32'ha135ee82;
    ram_cell[     634] = 32'hbc0e0347;
    ram_cell[     635] = 32'h9ac4a238;
    ram_cell[     636] = 32'hf00204de;
    ram_cell[     637] = 32'h2d56927e;
    ram_cell[     638] = 32'hd7404c66;
    ram_cell[     639] = 32'h2092408b;
    ram_cell[     640] = 32'h4268d370;
    ram_cell[     641] = 32'hfbe0c14c;
    ram_cell[     642] = 32'hdaa82d23;
    ram_cell[     643] = 32'hd5ebeee7;
    ram_cell[     644] = 32'h608563f8;
    ram_cell[     645] = 32'h16fe9812;
    ram_cell[     646] = 32'h63b26f75;
    ram_cell[     647] = 32'h8ac9fdcc;
    ram_cell[     648] = 32'h8d7d0ce7;
    ram_cell[     649] = 32'h22455125;
    ram_cell[     650] = 32'h844da6cd;
    ram_cell[     651] = 32'h63e6fe1b;
    ram_cell[     652] = 32'h1e4ffbaf;
    ram_cell[     653] = 32'had279841;
    ram_cell[     654] = 32'h86976411;
    ram_cell[     655] = 32'h57b78109;
    ram_cell[     656] = 32'hb66f1355;
    ram_cell[     657] = 32'hf9c68dee;
    ram_cell[     658] = 32'h0d829748;
    ram_cell[     659] = 32'ha8fed007;
    ram_cell[     660] = 32'h9aaec9c8;
    ram_cell[     661] = 32'h6d9932cd;
    ram_cell[     662] = 32'he4f4b94d;
    ram_cell[     663] = 32'h29d72aa6;
    ram_cell[     664] = 32'haef6b7fb;
    ram_cell[     665] = 32'hd2badf18;
    ram_cell[     666] = 32'h5c189160;
    ram_cell[     667] = 32'hfc103748;
    ram_cell[     668] = 32'hd5659231;
    ram_cell[     669] = 32'he32000fa;
    ram_cell[     670] = 32'h04e0999d;
    ram_cell[     671] = 32'h98d968e2;
    ram_cell[     672] = 32'h5567a1ca;
    ram_cell[     673] = 32'h8582a1f7;
    ram_cell[     674] = 32'hbb439384;
    ram_cell[     675] = 32'h966790ff;
    ram_cell[     676] = 32'h159e6664;
    ram_cell[     677] = 32'h66c826af;
    ram_cell[     678] = 32'h47afaa8e;
    ram_cell[     679] = 32'h3f602d12;
    ram_cell[     680] = 32'hbc1b5fa2;
    ram_cell[     681] = 32'h2e740bdc;
    ram_cell[     682] = 32'h9b5f1f5c;
    ram_cell[     683] = 32'ha3bb10d3;
    ram_cell[     684] = 32'h73aacf1d;
    ram_cell[     685] = 32'hcd2481bd;
    ram_cell[     686] = 32'hc0d44acf;
    ram_cell[     687] = 32'h548a9f03;
    ram_cell[     688] = 32'h5185b277;
    ram_cell[     689] = 32'h66c079f2;
    ram_cell[     690] = 32'h0a22cf6a;
    ram_cell[     691] = 32'h59fdf452;
    ram_cell[     692] = 32'hf7aa2711;
    ram_cell[     693] = 32'h529cdb8e;
    ram_cell[     694] = 32'h89517027;
    ram_cell[     695] = 32'h375f0122;
    ram_cell[     696] = 32'hce00fa7d;
    ram_cell[     697] = 32'hf0272dec;
    ram_cell[     698] = 32'h9d2c3f97;
    ram_cell[     699] = 32'h5b4ff6bb;
    ram_cell[     700] = 32'h2326dade;
    ram_cell[     701] = 32'hbc81514f;
    ram_cell[     702] = 32'h4e1c5a85;
    ram_cell[     703] = 32'h778b250b;
    ram_cell[     704] = 32'h534b85a1;
    ram_cell[     705] = 32'ha3df57d9;
    ram_cell[     706] = 32'h2164b4e5;
    ram_cell[     707] = 32'hba3f65e3;
    ram_cell[     708] = 32'hcd4985fa;
    ram_cell[     709] = 32'h64a23597;
    ram_cell[     710] = 32'h3e1aa411;
    ram_cell[     711] = 32'hf1ac8782;
    ram_cell[     712] = 32'hd5cc9bfd;
    ram_cell[     713] = 32'h5f40ffd4;
    ram_cell[     714] = 32'h57c85025;
    ram_cell[     715] = 32'h227d46ff;
    ram_cell[     716] = 32'h5045a252;
    ram_cell[     717] = 32'hb05f3f22;
    ram_cell[     718] = 32'h8b5c2b19;
    ram_cell[     719] = 32'hb77d636b;
    ram_cell[     720] = 32'h0ade71f7;
    ram_cell[     721] = 32'h8f338b3a;
    ram_cell[     722] = 32'hb1c060a4;
    ram_cell[     723] = 32'hbf1c12ed;
    ram_cell[     724] = 32'hf045f1b3;
    ram_cell[     725] = 32'hccd15b71;
    ram_cell[     726] = 32'h30156bca;
    ram_cell[     727] = 32'h4e8f7ec5;
    ram_cell[     728] = 32'h2176972b;
    ram_cell[     729] = 32'ha02fda90;
    ram_cell[     730] = 32'hc1416cee;
    ram_cell[     731] = 32'h4a6b064d;
    ram_cell[     732] = 32'h866c1f88;
    ram_cell[     733] = 32'h078bd6ca;
    ram_cell[     734] = 32'h9797c88a;
    ram_cell[     735] = 32'hf6f6855b;
    ram_cell[     736] = 32'h4637ea05;
    ram_cell[     737] = 32'h5788696d;
    ram_cell[     738] = 32'h42b237de;
    ram_cell[     739] = 32'h717bc602;
    ram_cell[     740] = 32'h6d2b1049;
    ram_cell[     741] = 32'h7be6b5a8;
    ram_cell[     742] = 32'hf7d80c45;
    ram_cell[     743] = 32'he747b456;
    ram_cell[     744] = 32'h7856acf8;
    ram_cell[     745] = 32'h470dc931;
    ram_cell[     746] = 32'h94baa6c7;
    ram_cell[     747] = 32'hdf0bbda9;
    ram_cell[     748] = 32'hfed20844;
    ram_cell[     749] = 32'h4a715150;
    ram_cell[     750] = 32'h439f2b9c;
    ram_cell[     751] = 32'h7609cdd3;
    ram_cell[     752] = 32'h9fb42574;
    ram_cell[     753] = 32'h4301a736;
    ram_cell[     754] = 32'h00904b41;
    ram_cell[     755] = 32'hc0f4608d;
    ram_cell[     756] = 32'h1442d579;
    ram_cell[     757] = 32'hd4975198;
    ram_cell[     758] = 32'h8555eb2a;
    ram_cell[     759] = 32'h94354fc6;
    ram_cell[     760] = 32'h2f14467d;
    ram_cell[     761] = 32'h54eaeb9a;
    ram_cell[     762] = 32'h09128f80;
    ram_cell[     763] = 32'h1ff60115;
    ram_cell[     764] = 32'hd5c350fb;
    ram_cell[     765] = 32'h4326ca42;
    ram_cell[     766] = 32'h096d9309;
    ram_cell[     767] = 32'hb223b2e9;
end

endmodule
